// +FHDR----------------------------------------------------------------------------
// Project Name  : Tiny RISC-V
// Author        : Qidc
// Email         : qidc@stu.pku.edu.cn
// Created On    : 2024/10/09 13:41
// Last Modified : 2024/10/09 13:41
// File Name     : inst_decode_tb.v
// Description   :
//         
// Copyright (c) 2024 Peking University.
// ALL RIGHTS RESERVED
// 
// ---------------------------------------------------------------------------------
// Modification History:
// Date         By              Version                 Change Description
// ---------------------------------------------------------------------------------
// 2024/10/09   Qidc            1.0                     Original
// -FHDR----------------------------------------------------------------------------
`timescale 1ns/1ps
module inst_decode_tb
(
);
endmodule

