// +FHDR----------------------------------------------------------------------------
// Project Name  : Tiny RISC-V
// Author        : Qidc
// Email         : qidc@stu.pku.edu.cn
// Created On    : 2024/10/09 13:39
// Last Modified : 2024/10/09 13:39
// File Name     : alu_tb.v
// Description   :
//         
// Copyright (c) 2024 Peking University.
// ALL RIGHTS RESERVED
// 
// ---------------------------------------------------------------------------------
// Modification History:
// Date         By              Version                 Change Description
// ---------------------------------------------------------------------------------
// 2024/10/09   Qidc            1.0                     Original
// -FHDR----------------------------------------------------------------------------
`timescale 1ns/1ps
module alu_tb
(
);
endmodule

